CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
220 200 30 200 9
1 79 853 1031
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
84 C:\Users\241pr\OneDrive - UBC\Desktop\UBC\ELEC 301\MP2\CircuitMaker60S\CM60S\BOM.DAT
0 7
1 79 853 1031
211550226 384
0
6 Title:
5 Name:
0
0
0
6
9 V Source~
197 540 378 0 2 5
0 3 2
0
0 0 17008 0
3 10V
13 0 34 8
3 Vce
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
8953 0 0
0
0
12 NPN Trans:B~
219 414 378 0 3 7
0 4 5 2
0
0 0 848 0
7 2N2222A
3 0 52 8
2 Q1
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 1 0 0
1 Q
4441 0 0
0
0
9 V Source~
197 279 387 0 2 5
0 6 2
0
0 0 17008 0
3 10V
13 -1 34 7
3 Vbe
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3618 0 0
0
0
7 Ground~
168 423 450 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
9 Resistor~
219 496 333 0 2 5
0 4 3
0
0 0 624 0
3 420
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 342 351 0 2 5
0 6 5
0
0 0 752 0
3 680
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
7
2 1 3 0 0 4224 0 5 1 0 0 3
514 333
540 333
540 357
1 1 4 0 0 8320 0 2 5 0 0 3
419 360
419 333
478 333
2 2 5 0 0 4224 0 6 2 0 0 4
360 351
388 351
388 378
396 378
1 1 6 0 0 8320 0 3 6 0 0 3
279 366
279 351
324 351
3 0 2 0 0 4096 0 2 0 0 6 3
419 396
419 410
423 410
1 2 2 0 0 8192 0 4 1 0 0 4
423 444
423 408
540 408
540 399
2 1 2 0 0 8320 0 3 4 0 0 4
279 408
279 436
423 436
423 444
0
0
2069 0 1
0
0
3 Vbe
0 0.7 0.01
3 Vce
0 10 0.01
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
4327268 1210432 100 100 0 0
0 0 0 0
1 79 162 149
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 5
0
1247232 8550464 100 100 0 0
77 66 797 396
853 79 1705 555
797 66
77 66
797 66
797 396
0 0
5e-006 0 5e-006 0 5e-006 5e-006
12385 0
4 1e-006 5
0
2427336 2259520 100 100 0 0
77 66 797 396
853 555 1705 1031
797 66
77 66
797 66
797 396
0 0
0.7 0 0.01 -0.002 0.7 0.7
12537 0
4 0.2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
