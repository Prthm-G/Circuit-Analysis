CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 200 30 200 9
0 71 2560 551
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
69 C:\Users\241pr\OneDrive - UBC\Desktop\Apps\UBC\ELEC 301\CM60S\BOM.DAT
0 7
0 71 2560 551
211288083 384
0
6 Title:
5 Name:
0
0
0
11
2 +V
167 452 413 0 1 3
0 8
0
0 0 53616 180
4 -15V
3 -7 31 1
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
2 +V
167 450 342 0 1 3
0 9
0
0 0 53616 0
3 15V
-7 -14 14 -6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
8 Op-Amp5~
219 450 378 0 5 11
0 2 5 9 8 6
0
0 0 80 0
5 UA741
43 -24 78 -16
2 U1
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 1 0 0
1 U
3618 0 0
0
0
10 Capacitor~
219 297 369 0 2 5
0 3 7
0
0 0 336 0
3 1uF
-11 -18 10 -10
1 C
-4 -28 3 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Capacitor~
219 207 369 0 2 5
0 4 3
0
0 0 848 0
3 1uF
-11 -18 10 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
10 Capacitor~
219 99 369 0 2 5
0 6 4
0
0 0 848 0
3 1uF
-11 -18 10 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
7 Ground~
168 396 450 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
9 Resistor~
219 450 306 0 2 5
0 5 6
0
0 0 880 0
5 29.1k
-17 -14 18 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 252 405 0 3 5
0 2 3 -1
0
0 0 368 90
2 1k
8 0 22 8
1 R
11 -10 18 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 144 405 0 3 5
0 2 4 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 369 369 0 2 5
0 7 5
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
14
2 0 3 0 0 4096 0 9 0 0 7 2
252 387
252 369
2 0 4 0 0 4096 0 10 0 0 6 2
144 387
144 369
1 0 5 0 0 8320 0 8 0 0 9 3
432 306
407 306
407 369
2 5 6 0 0 8192 0 8 3 0 0 4
468 306
476 306
476 378
468 378
1 2 6 0 0 12416 0 6 8 0 0 6
90 369
86 369
86 253
476 253
476 306
468 306
1 2 4 0 0 4224 0 5 6 0 0 2
198 369
108 369
1 2 3 0 0 4224 0 4 5 0 0 2
288 369
216 369
1 2 7 0 0 4224 0 11 4 0 0 2
351 369
306 369
2 2 5 0 0 0 0 11 3 0 0 4
387 369
424 369
424 372
432 372
1 0 2 0 0 8192 0 3 0 0 12 3
432 384
393 384
393 436
1 0 2 0 0 0 0 9 0 0 12 4
252 423
252 431
253 431
253 436
1 1 2 0 0 8320 0 10 7 0 0 4
144 423
144 436
396 436
396 444
4 1 8 0 0 4224 0 3 1 0 0 3
450 391
450 398
452 398
1 3 9 0 0 4224 0 2 3 0 0 2
450 351
450 365
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.1 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
853826 1210432 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 10
1
476 337
0 6 0 0 2	0 4 0 0
590570 8550976 100 100 0 0
77 66 2507 396
0 551 2560 1031
2507 66
77 66
2507 66
2507 396
0 0
0.1 0 0.00233218 0.00233206 0.1 0.1
12521 0
4 0.03 10
1
476 334
0 6 0 0 2	0 4 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
