CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
190 260 30 200 9
0 71 1024 1104
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
69 C:\Users\241pr\OneDrive - UBC\Desktop\Apps\UBC\ELEC 301\CM60S\BOM.DAT
0 7
0 71 1024 1104
211288083 384
0
6 Title:
5 Name:
0
0
0
22
7 Ground~
168 765 450 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
11 Signal Gen~
195 207 567 0 19 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1176256512 0 1020054733
20
1 10000 0 0.025 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -25m/25mV
-32 -30 31 -22
2 Vs
-7 -40 7 -32
0
0
39 %D %1 %2 DC 0 SIN(0 25m 10k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 360 459 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 252 612 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 702 612 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 612 612 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
10 Capacitor~
219 702 558 0 2 5
0 2 10
0
0 0 848 90
4 22uF
15 1 43 9
2 CE
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
10 Capacitor~
219 702 396 0 2 5
0 9 8
0
0 0 848 0
4 22uF
-14 -14 14 -6
3 CC2
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
10 Capacitor~
219 396 513 0 2 5
0 4 7
0
0 0 848 0
4 22uF
-15 -18 13 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
10 Capacitor~
219 396 423 0 2 5
0 2 6
0
0 0 848 0
5 150uF
-18 -18 17 -10
2 CB
-7 -31 7 -23
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7931 0 0
0
0
12 NPN Trans:B~
219 585 513 0 3 7
0 11 7 10
0
0 0 848 0
7 2N2222A
3 0 52 8
2 Q1
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 1 0 0
1 Q
9325 0 0
0
0
12 NPN Trans:B~
219 585 423 0 3 7
0 9 6 11
0
0 0 848 0
7 2N2222A
3 0 52 8
2 Q2
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 1 0 0
1 Q
8903 0 0
0
0
2 +V
167 531 333 0 1 3
0 12
0
0 0 54256 0
3 20V
-11 -22 10 -14
3 Vcc
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3834 0 0
0
0
7 Ground~
168 459 612 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
9 Resistor~
219 351 513 0 2 5
0 3 4
0
0 0 880 0
4 3.3k
-14 -15 14 -7
3 Rin
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 459 468 0 2 5
0 7 6
0
0 0 880 90
3 27k
5 0 26 8
3 RB2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 765 423 0 3 5
0 2 8 -1
0
0 0 880 90
3 50k
5 0 26 8
2 RL
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 297 513 0 2 5
0 5 3
0
0 0 880 0
2 50
-7 -14 7 -6
2 RS
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 612 558 0 3 5
0 2 10 -1
0
0 0 880 90
4 2.7k
1 0 29 8
2 RE
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 603 378 0 4 5
0 9 12 0 1
0
0 0 880 90
4 2.7k
1 0 29 8
2 RC
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 459 558 0 3 5
0 2 7 -1
0
0 0 880 90
3 36k
5 0 26 8
3 RB3
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 459 378 0 4 5
0 6 12 0 1
0
0 0 880 90
3 51k
5 1 26 9
3 RB1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
23
2 1 3 0 0 4224 0 18 15 0 0 2
315 513
333 513
2 1 4 0 0 4224 0 15 9 0 0 2
369 513
387 513
1 1 2 0 0 4096 0 17 1 0 0 2
765 441
765 444
2 1 2 0 0 8192 0 2 4 0 0 3
238 572
252 572
252 606
1 1 5 0 0 8320 0 2 18 0 0 4
238 562
252 562
252 513
279 513
1 1 2 0 0 0 0 3 10 0 0 3
360 453
360 423
387 423
2 0 6 0 0 4096 0 10 0 0 14 2
405 423
459 423
2 0 7 0 0 4096 0 9 0 0 13 2
405 513
460 513
2 2 8 0 0 8320 0 17 8 0 0 3
765 405
765 396
711 396
1 1 9 0 0 4224 0 8 20 0 0 5
693 396
611 396
611 404
603 404
603 396
1 1 2 0 0 4224 0 7 5 0 0 2
702 567
702 606
2 0 10 0 0 8320 0 7 0 0 16 3
702 549
702 535
612 535
2 0 7 0 0 4224 0 11 0 0 21 2
567 513
459 513
2 0 6 0 0 4224 0 12 0 0 22 2
567 423
459 423
1 1 2 0 0 0 0 19 6 0 0 2
612 576
612 606
3 2 10 0 0 0 0 11 19 0 0 4
590 531
590 535
612 535
612 540
3 1 11 0 0 8320 0 12 11 0 0 4
590 441
603 441
603 495
590 495
1 1 9 0 0 0 0 20 12 0 0 4
603 396
603 400
590 400
590 405
0 2 12 0 0 4224 0 0 20 23 0 3
531 352
603 352
603 360
1 1 2 0 0 0 0 21 14 0 0 2
459 576
459 606
1 2 7 0 0 0 0 16 21 0 0 2
459 486
459 540
1 2 6 0 0 0 0 22 16 0 0 2
459 396
459 450
1 2 12 0 0 0 0 13 22 0 0 4
531 342
531 352
459 352
459 360
0
0
2073 0 1
0
0
0
0 0 0
0
0 0 0
10 1 0.001 1e+011
0 0.0005 2e-006 2e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
656202 1210432 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 10
1
753 396
0 8 0 0 2	0 9 0 0
1182094 8550976 100 100 0 0
77 66 977 426
1024 71 2048 587
977 66
77 66
977 118
977 426
0 0
0.0005 0 4.26667e-006 -6e-006 0.0005 0.0005
12409 3
4 0.0001 10
0
1313238 4356162 100 100 0 0
77 66 987 426
1024 587 2048 1103
428 66
669 66
987 212
987 209
0 0
251.189 1.28142e+006 34 37 1e+011 1e+011
12530 0
4 3e+010 5e+010
1
756 396
0 8 0 0 2	0 9 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
