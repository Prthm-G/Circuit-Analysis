CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 10 30 200 9
1 79 853 1031
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
69 C:\Users\241pr\OneDrive - UBC\Desktop\Apps\UBC\ELEC 301\CM60S\BOM.DAT
0 7
1 79 853 1031
211288082 384
0
6 Title:
5 Name:
0
0
0
17
11 Signal Gen~
195 180 333 0 24 64
0 3 2 1 86 -10 10 9 0 0
0 0 0 0 0 0 0 1148846079 -1138501877 1008981771
0 814313567 814313567 973279855 981668463
20
0 1000 -0.01 0.01 0 1e-009 1e-009 0.0005 0.001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 336 0
9 -10m/10mV
-32 -30 31 -22
2 V3
-7 -40 7 -32
0
0
45 %D %1 %2 DC 0 PULSE(-10m 10m 0 1n 1n 500u 1m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
2 +V
167 424 59 0 1 3
0 12
0
0 0 53616 0
2 5V
-5 -15 9 -7
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
12 NPN Trans:B~
219 478 176 0 3 7
0 10 2 9
0
0 0 848 512
7 2N2222A
-57 0 -8 8
2 Q2
-39 -10 -25 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
3618 0 0
0
0
12 NPN Trans:B~
219 410 318 0 3 7
0 9 6 5
0
0 0 848 0
7 2N2222A
3 0 52 8
2 Q3
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
6153 0 0
0
0
12 NPN Trans:B~
219 364 177 0 3 7
0 11 8 9
0
0 0 848 0
7 2N2222A
3 0 52 8
2 Q4
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
5394 0 0
0
0
10 Capacitor~
219 334 320 0 2 5
0 7 6
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
7 Ground~
168 541 203 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
7 Ground~
168 325 248 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
7 Ground~
168 253 221 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3549 0 0
0
0
7 Ground~
168 235 365 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7931 0 0
0
0
2 +V
167 415 383 0 1 3
0 5
0
0 0 61680 180
3 -5V
6 -2 27 6
1 V
13 -12 20 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9325 0 0
0
0
11 Signal Gen~
195 190 194 0 64 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1203982336 0 1028443341
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -1338700788
20
1 100000 0 0.05 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 336 0
9 -50m/50mV
-32 -30 31 -22
2 V2
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 50m 100k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8903 0 0
0
0
9 Resistor~
219 370 113 0 4 5
0 11 12 0 1
0
0 0 368 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 469 113 0 4 5
0 10 12 0 1
0
0 0 368 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 307 176 0 2 5
0 4 8
0
0 0 368 0
2 50
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 370 266 0 4 5
0 6 2 0 -1
0
0 0 368 90
4 200k
1 0 29 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 271 320 0 2 5
0 3 7
0
0 0 368 0
2 2k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
17
2 1 2 0 0 4096 0 1 10 0 0 3
211 338
235 338
235 359
1 1 3 0 0 4224 0 1 17 0 0 4
211 328
245 328
245 320
253 320
2 1 2 0 0 4096 0 12 9 0 0 3
221 199
253 199
253 215
1 1 4 0 0 4224 0 12 15 0 0 4
221 189
281 189
281 176
289 176
1 3 5 0 0 4240 0 11 4 0 0 2
415 368
415 336
1 0 6 0 0 4112 0 16 0 0 9 2
370 284
370 320
1 2 2 0 0 8208 0 8 16 0 0 4
325 242
325 238
370 238
370 248
2 1 7 0 0 4240 0 17 6 0 0 2
289 320
325 320
2 2 6 0 0 4240 0 6 4 0 0 4
343 320
384 320
384 318
392 318
2 2 8 0 0 4240 0 5 15 0 0 4
346 177
333 177
333 176
325 176
0 1 9 0 0 4112 0 0 4 13 0 2
415 202
415 300
2 1 2 0 0 4240 0 3 7 0 0 3
492 176
541 176
541 197
3 3 9 0 0 8336 0 5 3 0 0 4
369 195
369 202
469 202
469 194
1 1 10 0 0 4240 0 14 3 0 0 2
469 131
469 158
1 1 11 0 0 4240 0 13 5 0 0 4
370 131
370 151
369 151
369 159
2 0 12 0 0 8208 0 14 0 0 17 3
469 95
469 87
424 87
1 2 12 0 0 8336 0 2 13 0 0 4
424 68
424 87
370 87
370 95
0
0
25 0 1
0
0
0
0 0 0
0
0 0 0
100 1 1 4e+009
0 0.5 1e-006 1e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1640056 1210432 100 100 0 0
0 0 0 0
1 79 162 149
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 3
0
3150312 8550976 5142 173 220 17
77 66 797 396
853 79 1705 555
797 66
797 66
797 66
797 66
469 147
0.231945 0.231945 3.65289 3.65289 0.5 0.5
12313 0
4 0.1 3
1
370 148
0 11 0 0 1	0 15 0 0
7669348 4356160 100 100 309 196
77 66 797 396
853 555 1705 1031
487 66
77 66
797 263
797 396
469 146
3.97554e+009 1.70854e+009 41.8727 24.9455 3.98107e+009 3.98107e+009
12401 0
4 1 20
1
370 144
0 11 0 0 1	0 15 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
