CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
360 200 30 200 9
0 71 1280 1032
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
69 C:\Users\241pr\OneDrive - UBC\Desktop\Apps\UBC\ELEC 301\CM60S\BOM.DAT
0 7
0 71 1280 1032
1285029907 384
0
6 Title:
5 Name:
0
0
0
29
5 SAVE-
218 878 580 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
22 *AC(dB) -1.000 1.000 0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
4 SAVE
8953 0 0
0
0
5 SAVE-
218 881 236 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
22 *AC(dB) -1.000 1.000 0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
4 SAVE
4441 0 0
0
0
10 Capacitor~
219 782 580 0 2 5
0 6 3
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C4
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
10 Capacitor~
219 440 580 0 2 5
0 4 5
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
2 +V
167 593 418 0 1 3
0 7
0
0 0 53616 0
3 15V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
7 Ground~
168 575 670 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
12 NPN Trans:B~
219 570 580 0 3 7
0 8 5 2
0
0 0 848 0
6 2N3904
7 1 49 9
2 Q4
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
9914 0 0
0
0
12 NPN Trans:B~
219 679 518 0 3 7
0 7 8 6
0
0 0 848 0
6 2N3904
7 0 49 8
2 Q3
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
3747 0 0
0
0
11 Signal Gen~
195 242 634 0 64 64
0 9 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 981668463
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 106026014
20
1 1000 0 0.001 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -1m/1mV
-25 -30 24 -22
2 V3
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
11 Signal Gen~
195 242 290 0 64 64
0 16 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 981668463
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 106026014
20
1 1000 0 0.001 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -1m/1mV
-25 -30 24 -22
2 V1
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
12 NPN Trans:B~
219 679 174 0 3 7
0 14 15 13
0
0 0 848 0
6 2N3904
7 0 49 8
2 Q2
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
9325 0 0
0
0
12 NPN Trans:B~
219 570 236 0 3 7
0 15 12 2
0
0 0 848 0
6 2N3904
7 1 49 9
2 Q1
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
8903 0 0
0
0
7 Ground~
168 575 326 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
2 +V
167 593 74 0 1 3
0 14
0
0 0 53616 0
3 15V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
10 Capacitor~
219 440 236 0 2 5
0 11 12
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7668 0 0
0
0
10 Capacitor~
219 782 236 0 2 5
0 13 10
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4718 0 0
0
0
9 Resistor~
219 593 733 0 2 5
0 4 3
0
0 0 752 0
4 100k
-15 -14 13 -6
3 Rf1
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 908 616 0 3 5
0 2 3 -1
0
0 0 880 90
3 10k
5 0 26 8
3 RL1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 485 625 0 3 5
0 2 5 -1
0
0 0 880 90
3 20k
5 -2 26 6
3 RB1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 683 625 0 3 5
0 2 6 -1
0
0 0 880 90
3 560
8 0 29 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 593 472 0 4 5
0 8 7 0 1
0
0 0 880 90
3 10k
5 0 26 8
3 Rc1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 485 472 0 4 5
0 5 7 0 1
0
0 0 880 90
4 330k
1 0 29 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 350 580 0 2 5
0 9 4
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 350 236 0 2 5
0 16 11
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 485 128 0 4 5
0 12 14 0 1
0
0 0 880 90
4 330k
1 0 29 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
9 Resistor~
219 593 128 0 4 5
0 15 14 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 Rc
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
9 Resistor~
219 683 281 0 3 5
0 2 13 -1
0
0 0 880 90
3 560
8 0 29 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5670 0 0
0
0
9 Resistor~
219 485 281 0 3 5
0 2 12 -1
0
0 0 880 90
3 20k
5 -2 26 6
3 RB2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 908 272 0 3 5
0 2 10 -1
0
0 0 880 90
3 10k
5 0 26 8
2 RL
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
42
1 0 2 0 0 4096 0 20 0 0 14 2
683 643
683 655
0 0 2 0 0 4096 0 0 0 12 16 2
485 654
575 654
2 0 3 0 0 4224 0 17 0 0 8 3
611 733
856 733
856 580
0 1 4 0 0 8320 0 0 17 10 0 3
386 580
386 733
575 733
2 0 5 0 0 4096 0 19 0 0 6 3
485 607
485 579
486 579
1 0 5 0 0 4096 0 22 0 0 7 4
485 490
485 575
486 575
486 580
2 2 5 0 0 4224 0 4 7 0 0 2
449 580
552 580
2 2 3 0 0 0 0 3 18 0 0 3
791 580
908 580
908 598
0 1 6 0 0 4224 0 0 3 15 0 2
684 580
773 580
2 1 4 0 0 0 0 23 4 0 0 2
368 580
431 580
1 0 7 0 0 4096 0 5 0 0 19 2
593 427
593 445
1 2 2 0 0 16384 0 19 9 0 0 5
485 643
485 664
477 664
477 639
273 639
1 0 2 0 0 0 0 6 0 0 16 2
575 664
575 664
1 0 2 0 0 8320 0 18 0 0 16 3
908 634
908 655
575 655
2 3 6 0 0 0 0 20 8 0 0 3
683 607
684 607
684 536
3 0 2 0 0 0 0 7 0 0 0 2
575 598
575 670
0 2 8 0 0 4096 0 0 8 18 0 2
592 518
661 518
1 1 8 0 0 8320 0 7 21 0 0 4
575 562
592 562
592 490
593 490
0 1 7 0 0 8192 0 0 8 20 0 4
593 446
593 445
684 445
684 500
2 2 7 0 0 8320 0 22 21 0 0 4
485 454
485 446
593 446
593 454
1 1 9 0 0 4224 0 9 23 0 0 4
273 629
324 629
324 580
332 580
1 0 2 0 0 0 0 27 0 0 35 2
683 299
683 311
0 0 2 0 0 0 0 0 0 33 37 2
485 310
575 310
0 0 10 0 0 4224 0 0 0 0 29 3
611 389
856 389
856 236
0 0 11 0 0 8320 0 0 0 31 0 3
386 236
386 389
575 389
2 0 12 0 0 4096 0 28 0 0 27 3
485 263
485 235
486 235
1 0 12 0 0 4096 0 25 0 0 28 4
485 146
485 231
486 231
486 236
2 2 12 0 0 4224 0 15 12 0 0 2
449 236
552 236
2 2 10 0 0 0 0 16 29 0 0 3
791 236
908 236
908 254
0 1 13 0 0 4224 0 0 16 36 0 2
684 236
773 236
2 1 11 0 0 0 0 24 15 0 0 2
368 236
431 236
1 0 14 0 0 4096 0 14 0 0 40 2
593 83
593 101
1 2 2 0 0 0 0 28 10 0 0 5
485 299
485 320
477 320
477 295
273 295
1 0 2 0 0 0 0 13 0 0 37 2
575 320
575 320
1 0 2 0 0 0 0 29 0 0 37 3
908 290
908 311
575 311
2 3 13 0 0 0 0 27 11 0 0 3
683 263
684 263
684 192
3 0 2 0 0 0 0 12 0 0 0 2
575 254
575 326
0 2 15 0 0 4096 0 0 11 39 0 2
592 174
661 174
1 1 15 0 0 8320 0 12 26 0 0 4
575 218
592 218
592 146
593 146
0 1 14 0 0 8192 0 0 11 41 0 4
593 102
593 101
684 101
684 156
2 2 14 0 0 8320 0 25 26 0 0 4
485 110
485 102
593 102
593 110
1 1 16 0 0 4224 0 10 24 0 0 4
273 285
324 285
324 236
332 236
0
0
2073 0 1
0
0
0
0 0 0
0
0 0 0
100 1 0.01 1e+008
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
2 0 0 0
2 Rc
9900 10100 100
3 Rc1
9900 10100 100
5 -1 10 10 10 0 10 10 0
8325386 1079360 100 100 0 0
0 0 0 0
422 84 583 154
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 10
0
11405712 8813120 100 100 0 0
77 66 1247 396
1280 71 2560 551
1247 66
77 66
1247 66
1247 396
0 0
0.005 0 0.005 0 0.005 0.005
28921 0
4 0.001 10
0
14158116 4290624 9999 2892 1011 557
77 66 2527 876
0 71 2560 1032
77 66
77 66
2527 66
2527 444
0 0
0.628148 0.628148 41.8182 24.7333 1e+008 1e+008
12530 0
4 3e+007 5e+007
20
856 598
0 3 0 0 2	0 3 0 0
856 598
0 3 0 0 2	0 3 0 0
856 598
0 3 0 0 2	0 3 0 0
856 598
0 3 0 0 2	0 3 0 0
856 598
0 3 0 0 2	0 3 0 0
856 598
0 3 0 0 2	0 3 0 0
856 598
0 3 0 0 2	0 3 0 0
856 598
0 3 0 0 2	0 3 0 0
856 598
0 3 0 0 2	0 3 0 0
856 598
0 3 0 0 2	0 3 0 0
882 236
0 10 0 0 1	0 29 0 0
882 236
0 10 0 0 1	0 29 0 0
882 236
0 10 0 0 1	0 29 0 0
882 236
0 10 0 0 1	0 29 0 0
882 236
0 10 0 0 1	0 29 0 0
882 236
0 10 0 0 1	0 29 0 0
882 236
0 10 0 0 1	0 29 0 0
882 236
0 10 0 0 1	0 29 0 0
882 236
0 10 0 0 1	0 29 0 0
882 236
0 10 0 0 1	0 29 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
