CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
230 180 30 200 9
1281 79 2133 1031
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
69 C:\Users\241pr\OneDrive - UBC\Desktop\Apps\UBC\ELEC 301\CM60S\BOM.DAT
0 7
1281 79 2133 1031
211288082 384
0
6 Title:
5 Name:
0
0
0
12
7 Ground~
168 324 414 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
2 +V
167 549 405 0 1 3
0 3
0
0 0 53616 180
3 -15
8 -18 29 -10
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
2 +V
167 549 324 0 1 3
0 4
0
0 0 53616 0
3 +15
-28 0 -7 8
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3618 0 0
0
0
7 Ground~
168 405 297 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
8 Op-Amp5~
219 549 360 0 5 11
0 7 6 4 3 5
0
0 0 848 0
5 UA741
19 -25 54 -17
2 U1
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 1 0 0
1 U
5394 0 0
0
0
10 Capacitor~
219 486 414 0 2 5
0 2 7
0
0 0 848 90
5 1.6nF
12 0 47 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
10 Capacitor~
219 396 414 0 2 5
0 5 8
0
0 0 848 90
5 1.6nF
11 0 46 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
7 Ground~
168 486 450 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
9 Resistor~
219 540 279 0 2 5
0 6 5
0
0 0 880 0
6 6.667k
-21 -14 21 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 432 279 0 3 5
0 2 6 -1
0
0 0 880 0
6 3.333k
-21 -14 21 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 432 369 0 2 5
0 8 7
0
0 0 368 0
3 10k
-10 -14 11 -6
1 R
-4 -24 3 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 351 369 0 3 5
0 2 8 -1
0
0 0 368 0
3 10k
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
13
1 1 2 0 0 4224 0 1 12 0 0 3
324 408
324 369
333 369
1 4 3 0 0 4224 0 2 5 0 0 2
549 390
549 373
1 3 4 0 0 4224 0 3 5 0 0 2
549 333
549 347
2 0 5 0 0 8192 0 9 0 0 11 3
558 279
611 279
611 360
2 0 6 0 0 8320 0 5 0 0 9 3
531 354
486 354
486 279
1 1 2 0 0 128 0 6 8 0 0 2
486 423
486 444
2 0 7 0 0 4096 0 6 0 0 8 2
486 405
486 369
2 1 7 0 0 4224 0 11 5 0 0 3
450 369
531 369
531 366
2 1 6 0 0 0 0 10 9 0 0 2
450 279
522 279
1 1 2 0 0 0 0 4 10 0 0 3
405 291
405 279
414 279
1 5 5 0 0 8320 0 7 5 0 0 5
396 423
396 495
611 495
611 360
567 360
2 0 8 0 0 4096 0 7 0 0 13 2
396 405
396 369
2 1 8 0 0 4224 0 12 11 0 0 2
369 369
414 369
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
100 1 1 1e+009
0 0.001 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
24250776 1210432 100 100 0 0
0 0 0 0
693 83 854 153
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 10
0
5703350 8550976 100 100 0 0
77 66 1667 876
1281 79 2986 1031
1617 66
119 66
1667 101
1667 847
0 0
0.000968917 2.68755e-005 -0.00421905 -0.00421911 0.001 0.001
12537 1
4 0.001 10
1
606 360
0 5 0 0 4	0 11 0 0
4655376 4421696 100 100 0 0
77 66 815 396
854 563 1706 1039
810 66
77 66
815 122
815 73
0 0
8.69009e+008 1 -0.0363636 8 1e+009 1e+009
12530 0
4 3e+011 5e+011
1
611 360
0 6 0 0 2	0 4 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
