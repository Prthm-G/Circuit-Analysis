CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
140 260 30 200 9
1 79 853 1031
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
69 C:\Users\241pr\OneDrive - UBC\Desktop\Apps\UBC\ELEC 301\CM60S\BOM.DAT
0 7
1 79 853 1031
211288082 384
0
6 Title:
5 Name:
0
0
0
14
7 Ground~
168 576 441 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 243 450 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 288 504 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
2 +V
167 369 666 0 1 3
0 5
0
0 0 53616 180
4 -12V
-13 2 15 10
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
12 NPN Trans:B~
219 423 603 0 3 7
0 7 6 5
0
0 0 848 0
7 2N2222A
3 0 52 8
2 Q4
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
5394 0 0
0
0
12 NPN Trans:B~
219 324 603 0 3 7
0 6 6 5
0
0 0 848 512
7 2N2222A
-57 0 -8 8
2 Q3
-39 -10 -25 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
7734 0 0
0
0
2 +V
167 441 252 0 1 3
0 3
0
0 0 53616 0
3 12V
-9 -15 12 -7
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
12 NPN Trans:B~
219 513 396 0 3 7
0 4 2 7
0
0 0 848 512
7 2N2222A
-57 0 -8 8
2 Q2
-39 -10 -25 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
3747 0 0
0
0
12 NPN Trans:B~
219 369 396 0 3 7
0 8 9 7
0
0 0 848 0
7 2N2222A
17 0 66 8
2 Q1
35 -10 49 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
3549 0 0
0
0
11 Signal Gen~
195 189 423 0 19 64
0 10 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1203982336 0 1050253722
20
1 100000 0 0.3 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 336 0
11 -300m/300mV
-39 -30 38 -22
2 V1
-7 -40 7 -32
0
0
41 %D %1 %2 DC 0 SIN(0 300m 100k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
9 Resistor~
219 315 531 0 4 5
0 6 2 0 -1
0
0 0 368 90
4 5.6k
2 0 30 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 504 315 0 4 5
0 4 3 0 1
0
0 0 368 90
2 8k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 378 315 0 4 5
0 8 3 0 1
0
0 0 368 90
2 8k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 297 396 0 2 5
0 10 9
0
0 0 368 0
2 50
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
16
2 1 2 0 0 4224 0 8 1 0 0 3
527 396
576 396
576 435
2 1 2 0 0 0 0 10 2 0 0 3
220 428
243 428
243 444
1 0 3 0 0 4096 0 7 0 0 4 2
441 261
441 289
2 2 3 0 0 8320 0 13 12 0 0 4
378 297
378 289
504 289
504 297
1 1 4 0 0 4224 0 12 8 0 0 2
504 333
504 378
1 0 5 0 0 4096 0 4 0 0 10 2
369 651
369 629
0 0 6 0 0 4096 0 0 0 9 8 3
315 568
371 568
371 603
2 2 6 0 0 4224 0 6 5 0 0 2
338 603
405 603
1 1 6 0 0 0 0 11 6 0 0 2
315 549
315 585
3 3 5 0 0 8320 0 6 5 0 0 4
315 621
315 629
428 629
428 621
1 0 7 0 0 4224 0 5 0 0 12 2
428 585
428 422
3 3 7 0 0 0 0 9 8 0 0 4
374 414
374 422
504 422
504 414
1 1 8 0 0 4224 0 9 13 0 0 4
374 378
374 341
378 341
378 333
2 2 9 0 0 4224 0 14 9 0 0 2
315 396
351 396
1 1 10 0 0 4224 0 10 14 0 0 4
220 418
271 418
271 396
279 396
1 2 2 0 0 0 0 3 11 0 0 3
288 512
288 513
315 513
0
0
2065 0 2
0
0
0
0 0 0
0
0 0 0
100 1 1 1e+010
0 5e-005 2e-007 2e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
8983508 1210432 100 100 0 0
0 0 0 0
1 84 162 154
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 5
1
261 418
0 10 0 0 1	0 15 0 0
11797960 8550464 100 100 0 0
77 66 797 396
853 79 1705 555
797 66
77 66
797 178
797 345
504 345
5e-005 0 0.0963636 -0.207273 5e-005 5e-005
12401 0
4 0.001 5
1
255 418
0 10 0 0 1	0 15 0 0
20188494 4421696 355 523 318 196
77 66 817 396
853 555 1705 1031
770 66
770 66
817 219
817 262
0 0
8.55919e+006 8.55919e+006 43.6489 40.6591 1e+010 1e+010
12530 0
4 3e+009 5e+009
1
374 356
0 8 0 0 1	0 13 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
