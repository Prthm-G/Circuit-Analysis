CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
240 200 30 200 9
918 114 3350 1005
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
84 C:\Users\241pr\OneDrive - UBC\Desktop\UBC\ELEC 301\MP2\CircuitMaker60S\CM60S\BOM.DAT
0 7
918 114 3350 1005
211288082 384
0
6 Title:
5 Name:
0
0
0
5
9 V Source~
197 495 432 0 2 5
0 3 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
8953 0 0
0
0
9 V Source~
197 315 432 0 2 5
0 5 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
4441 0 0
0
0
12 NPN Trans:B~
219 378 396 0 3 7
0 4 5 2
0
0 0 848 0
7 2N2222A
3 0 52 8
2 Q1
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
3618 0 0
0
0
7 Ground~
168 414 459 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
9 Resistor~
219 450 342 0 2 5
0 4 3
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
6
3 0 2 0 0 4096 0 3 0 0 2 3
383 414
383 449
414 449
1 2 2 0 0 8192 0 4 1 0 0 6
414 453
414 449
481 449
481 459
495 459
495 453
2 1 2 0 0 8320 0 2 4 0 0 6
315 453
315 458
401 458
401 448
414 448
414 453
2 1 3 0 0 8320 0 5 1 0 0 3
468 342
495 342
495 411
1 1 4 0 0 8320 0 3 5 0 0 3
383 378
383 342
432 342
1 2 5 0 0 8320 0 2 3 0 0 3
315 411
315 396
360 396
0
0
2069 0 1
0
0
3 Vs1
0 3 0.02
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
