CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
180 140 30 200 9
0 71 2048 1104
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
69 C:\Users\241pr\OneDrive - UBC\Desktop\Apps\UBC\ELEC 301\CM60S\BOM.DAT
0 7
0 71 2048 1104
211288082 384
0
6 Title:
5 Name:
0
0
0
17
7 Ground~
168 1053 432 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
11 Signal Gen~
195 486 369 0 19 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1203982336 0 981668463
20
1 100000 0 0.001 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -1m/1mV
-25 -30 24 -22
2 V1
-7 -40 7 -32
0
0
39 %D %1 %2 DC 0 SIN(0 1m 100k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 927 432 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
2 +V
167 927 171 0 1 3
0 7
0
0 0 54256 0
3 12V
-11 -22 10 -14
3 Vcc
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
7 Ground~
168 594 207 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
10 Capacitor~
219 981 351 0 2 5
0 5 3
0
0 0 848 0
5 4.7uF
-18 -18 17 -10
3 Cc2
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
12 NPN Trans:B~
219 918 315 0 3 7
0 7 6 5
0
0 0 848 0
6 2N3904
7 0 49 8
2 Q2
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
9914 0 0
0
0
12 NPN Trans:B~
219 684 306 0 3 7
0 6 8 9
0
0 0 848 270
6 2N3904
-23 30 19 38
2 Q1
-9 20 5 28
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3747 0 0
0
0
10 Capacitor~
219 756 243 0 2 5
0 8 2
0
0 0 848 90
7 0.082uF
4 11 53 19
2 CB
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
10 Capacitor~
219 585 315 0 2 5
0 4 9
0
0 0 848 0
5 4.7uF
-19 -18 16 -10
3 Cc1
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7931 0 0
0
0
7 Ground~
168 531 432 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
9 Resistor~
219 1053 378 0 3 5
0 2 3 -1
0
0 0 880 90
2 50
8 0 22 8
2 RL
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 927 387 0 3 5
0 2 5 -1
0
0 0 880 90
4 1.6k
1 0 29 8
3 RE2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 873 243 0 4 5
0 6 7 0 1
0
0 0 880 90
4 7.5k
1 0 29 8
3 RC1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 819 243 0 4 5
0 8 7 0 1
0
0 0 880 90
4 150k
1 0 29 8
3 RB1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 684 243 0 4 5
0 8 2 0 -1
0
0 0 880 90
4 100k
1 0 29 8
3 RB2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 630 243 0 4 5
0 9 2 0 -1
0
0 0 880 90
4 7.5k
1 0 29 8
3 RE1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
20
1 1 2 0 0 4096 0 12 1 0 0 2
1053 396
1053 426
2 2 3 0 0 4224 0 6 12 0 0 3
990 351
1053 351
1053 360
1 1 4 0 0 4224 0 2 10 0 0 4
517 364
568 364
568 315
576 315
1 1 2 0 0 0 0 13 3 0 0 2
927 405
927 426
2 0 5 0 0 4096 0 13 0 0 18 4
927 369
927 356
928 356
928 351
1 0 6 0 0 4096 0 14 0 0 8 2
873 261
873 313
0 1 7 0 0 4224 0 0 7 10 0 2
923 188
923 297
1 2 6 0 0 4224 0 8 7 0 0 4
700 313
892 313
892 315
900 315
2 0 7 0 0 0 0 14 0 0 10 2
873 225
873 188
2 1 7 0 0 0 0 15 4 0 0 4
819 225
819 188
927 188
927 180
0 1 8 0 0 4096 0 0 15 17 0 3
756 282
819 282
819 261
2 0 2 0 0 0 0 16 0 0 14 4
684 225
684 198
685 198
685 193
2 0 2 0 0 0 0 17 0 0 14 4
630 225
630 198
631 198
631 193
2 1 2 0 0 8320 0 9 5 0 0 4
756 234
756 193
594 193
594 201
1 0 9 0 0 4096 0 17 0 0 19 2
630 261
630 315
1 0 8 0 0 0 0 16 0 0 17 2
684 261
684 282
1 2 8 0 0 8320 0 9 8 0 0 4
756 252
756 282
682 282
682 290
3 1 5 0 0 8320 0 7 6 0 0 3
923 333
923 351
972 351
2 3 9 0 0 4224 0 10 8 0 0 4
594 315
656 315
656 313
664 313
2 1 2 0 0 0 0 2 11 0 0 5
517 374
526 374
526 390
531 390
531 426
0
0
2065 0 2
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-005 2e-007 2e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
28380890 1079360 100 100 0 0
0 0 0 0
51 145 212 215
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 10
1
559 364
0 4 0 0 1	0 3 0 0
13112076 8550464 100 100 0 0
77 66 1997 936
0 71 2048 1104
1997 66
77 66
1997 91
1997 936
504 355
5e-005 0 1.98414e-005 -2.1e-005 5e-005 5e-005
12401 3
4 1e-005 10
0
5116706 4421696 100 100 0 0
77 66 1672 876
1 79 1706 1031
512 66
1027 66
1672 93
1672 114
0 0
8.64842e+006 8.64842e+006 43.6946 40.692 1e+010 1e+010
12530 0
4 3e+010 5e+010
1
1051 351
0 3 0 0 1	0 2 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
