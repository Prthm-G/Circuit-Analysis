CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
690 320 30 250 9
1 79 1025 1112
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
69 C:\Users\241pr\OneDrive - UBC\Desktop\Apps\UBC\ELEC 301\CM60S\BOM.DAT
0 7
1 79 1025 1112
1285029906 384
0
6 Title:
5 Name:
0
0
0
44
11 Signal Gen~
195 174 1026 0 64 64
0 9 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 981668463
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -1355074619
20
1 1000 0 0.001 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -1m/1mV
-25 -30 24 -22
2 V6
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
12 NPN Trans:B~
219 611 910 0 3 7
0 7 8 6
0
0 0 848 0
6 2N3904
7 0 49 8
2 Q6
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
4441 0 0
0
0
12 NPN Trans:B~
219 502 972 0 3 7
0 8 5 2
0
0 0 848 0
6 2N3904
7 1 49 9
2 Q5
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
3618 0 0
0
0
7 Ground~
168 507 1062 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
2 +V
167 525 810 0 1 3
0 7
0
0 0 53616 0
3 15V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
10 Capacitor~
219 372 972 0 2 5
0 4 5
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C6
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
10 Capacitor~
219 714 972 0 2 5
0 6 3
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C5
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
11 Signal Gen~
195 167 679 0 64 64
0 16 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 981668463
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -2009386014
20
1 1000 0 0.001 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -1m/1mV
-25 -30 24 -22
2 V4
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
12 NPN Trans:B~
219 604 563 0 3 7
0 14 15 13
0
0 0 848 0
6 2N3904
7 0 49 8
2 Q4
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
3549 0 0
0
0
12 NPN Trans:B~
219 495 625 0 3 7
0 15 12 2
0
0 0 848 0
6 2N3904
7 1 49 9
2 Q3
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
7931 0 0
0
0
7 Ground~
168 500 715 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
2 +V
167 518 463 0 1 3
0 14
0
0 0 53616 0
3 15V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
10 Capacitor~
219 365 625 0 2 5
0 11 12
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C4
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3834 0 0
0
0
10 Capacitor~
219 707 625 0 2 5
0 13 10
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3363 0 0
0
0
5 SAVE-
218 795 625 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
22 *AC(dB) -1.000 1.000 0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
7668 0 0
0
0
5 SAVE-
218 799 270 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
22 *AC(dB) -1.000 1.000 0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
4718 0 0
0
0
10 Capacitor~
219 711 270 0 2 5
0 20 17
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3874 0 0
0
0
10 Capacitor~
219 369 270 0 2 5
0 18 19
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6671 0 0
0
0
2 +V
167 522 108 0 1 3
0 21
0
0 0 53616 0
3 15V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3789 0 0
0
0
7 Ground~
168 504 360 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4871 0 0
0
0
12 NPN Trans:B~
219 499 270 0 3 7
0 22 19 2
0
0 0 848 0
6 2N3904
7 1 49 9
2 Q1
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
3750 0 0
0
0
12 NPN Trans:B~
219 608 208 0 3 7
0 21 22 20
0
0 0 848 0
6 2N3904
7 0 49 8
2 Q2
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
8778 0 0
0
0
11 Signal Gen~
195 171 324 0 19 64
0 23 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 981668463
20
1 1000 0 0.001 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -1m/1mV
-25 -30 24 -22
2 V1
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
538 0 0
0
0
9 Resistor~
219 282 972 0 2 5
0 9 4
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 417 864 0 4 5
0 5 7 0 1
0
0 0 880 90
4 330k
1 0 29 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
9 Resistor~
219 525 864 0 4 5
0 8 7 0 1
0
0 0 880 90
3 10k
5 0 26 8
3 Rc2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
9 Resistor~
219 615 1017 0 3 5
0 2 6 -1
0
0 0 880 90
3 560
8 0 29 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5670 0 0
0
0
9 Resistor~
219 417 1017 0 3 5
0 2 5 -1
0
0 0 880 90
3 20k
5 -2 26 6
3 RB3
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 840 1008 0 3 5
0 2 3 -1
0
0 0 880 90
3 10k
5 0 26 8
3 RL2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 525 1125 0 2 5
0 4 3
0
0 0 752 0
4 100k
-15 -14 13 -6
3 Rf2
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 275 625 0 2 5
0 16 11
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 410 517 0 4 5
0 12 14 0 1
0
0 0 880 90
4 330k
1 0 29 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
9 Resistor~
219 518 517 0 4 5
0 15 14 0 1
0
0 0 880 90
3 10k
5 0 26 8
3 Rc1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3635 0 0
0
0
9 Resistor~
219 608 670 0 3 5
0 2 13 -1
0
0 0 880 90
3 560
8 0 29 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3973 0 0
0
0
9 Resistor~
219 410 670 0 3 5
0 2 12 -1
0
0 0 880 90
3 20k
5 -2 26 6
3 RB1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
3851 0 0
0
0
9 Resistor~
219 833 661 0 3 5
0 2 10 -1
0
0 0 880 90
3 10k
5 0 26 8
3 RL1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8383 0 0
0
0
9 Resistor~
219 518 778 0 2 5
0 11 10
0
0 0 752 0
2 1k
-8 -14 6 -6
3 Rf1
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
9 Resistor~
219 522 423 0 2 5
0 18 17
0
0 0 752 0
2 1k
-8 -14 6 -6
2 Rf
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 837 306 0 3 5
0 2 17 -1
0
0 0 880 90
3 10k
5 0 26 8
2 RL
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3334 0 0
0
0
9 Resistor~
219 414 315 0 3 5
0 2 19 -1
0
0 0 880 90
3 20k
5 -2 26 6
3 RB2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
3559 0 0
0
0
9 Resistor~
219 612 315 0 3 5
0 2 20 -1
0
0 0 880 90
3 560
8 0 29 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
984 0 0
0
0
9 Resistor~
219 522 162 0 4 5
0 22 21 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 Rc
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7557 0 0
0
0
9 Resistor~
219 414 162 0 4 5
0 19 21 0 1
0
0 0 880 90
4 330k
1 0 29 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3146 0 0
0
0
9 Resistor~
219 279 270 0 2 5
0 23 18
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5687 0 0
0
0
63
1 0 2 0 0 4112 0 27 0 0 14 2
615 1035
615 1047
0 0 2 0 0 4112 0 0 0 12 16 2
417 1046
507 1046
2 0 3 0 0 4240 0 30 0 0 8 3
543 1125
788 1125
788 972
0 1 4 0 0 8336 0 0 30 10 0 3
318 972
318 1125
507 1125
2 0 5 0 0 4112 0 28 0 0 6 3
417 999
417 971
418 971
1 0 5 0 0 4112 0 25 0 0 7 4
417 882
417 967
418 967
418 972
2 2 5 0 0 4240 0 6 3 0 0 2
381 972
484 972
2 2 3 0 0 16 0 7 29 0 0 3
723 972
840 972
840 990
0 1 6 0 0 4240 0 0 7 15 0 2
616 972
705 972
2 1 4 0 0 16 0 24 6 0 0 2
300 972
363 972
1 0 7 0 0 4112 0 5 0 0 19 2
525 819
525 837
1 2 2 0 0 16400 0 28 1 0 0 5
417 1035
417 1056
409 1056
409 1031
205 1031
1 0 2 0 0 16 0 4 0 0 16 2
507 1056
507 1056
1 0 2 0 0 8336 0 29 0 0 16 3
840 1026
840 1047
507 1047
2 3 6 0 0 16 0 27 2 0 0 3
615 999
616 999
616 928
3 0 2 0 0 16 0 3 0 0 0 2
507 990
507 1062
0 2 8 0 0 4112 0 0 2 18 0 2
524 910
593 910
1 1 8 0 0 8336 0 3 26 0 0 4
507 954
524 954
524 882
525 882
0 1 7 0 0 8208 0 0 2 20 0 4
525 838
525 837
616 837
616 892
2 2 7 0 0 8336 0 25 26 0 0 4
417 846
417 838
525 838
525 846
1 1 9 0 0 4240 0 1 24 0 0 4
205 1021
256 1021
256 972
264 972
1 0 2 0 0 0 0 34 0 0 35 2
608 688
608 700
0 0 2 0 0 0 0 0 0 33 37 2
410 699
500 699
2 0 10 0 0 4224 0 37 0 0 29 3
536 778
781 778
781 625
0 1 11 0 0 8320 0 0 37 31 0 3
311 625
311 778
500 778
2 0 12 0 0 4096 0 35 0 0 27 3
410 652
410 624
411 624
1 0 12 0 0 4096 0 32 0 0 28 4
410 535
410 620
411 620
411 625
2 2 12 0 0 4224 0 13 10 0 0 2
374 625
477 625
2 2 10 0 0 0 0 14 36 0 0 3
716 625
833 625
833 643
0 1 13 0 0 4224 0 0 14 36 0 2
609 625
698 625
2 1 11 0 0 0 0 31 13 0 0 2
293 625
356 625
1 0 14 0 0 4096 0 12 0 0 40 2
518 472
518 490
1 2 2 0 0 0 0 35 8 0 0 5
410 688
410 709
402 709
402 684
198 684
1 0 2 0 0 0 0 11 0 0 37 2
500 709
500 709
1 0 2 0 0 0 0 36 0 0 37 3
833 679
833 700
500 700
2 3 13 0 0 0 0 34 9 0 0 3
608 652
609 652
609 581
3 0 2 0 0 0 0 10 0 0 0 2
500 643
500 715
0 2 15 0 0 4096 0 0 9 39 0 2
517 563
586 563
1 1 15 0 0 8320 0 10 33 0 0 4
500 607
517 607
517 535
518 535
0 1 14 0 0 8192 0 0 9 41 0 4
518 491
518 490
609 490
609 545
2 2 14 0 0 8320 0 32 33 0 0 4
410 499
410 491
518 491
518 499
1 1 16 0 0 4224 0 8 31 0 0 4
198 674
249 674
249 625
257 625
1 0 2 0 0 0 0 41 0 0 56 2
612 333
612 345
0 0 2 0 0 0 0 0 0 54 58 2
414 344
504 344
2 0 17 0 0 4224 0 38 0 0 50 3
540 423
785 423
785 270
0 1 18 0 0 8320 0 0 38 52 0 3
315 270
315 423
504 423
2 0 19 0 0 4096 0 40 0 0 48 3
414 297
414 269
415 269
1 0 19 0 0 4096 0 43 0 0 49 4
414 180
414 265
415 265
415 270
2 2 19 0 0 4224 0 18 21 0 0 2
378 270
481 270
2 2 17 0 0 0 0 17 39 0 0 3
720 270
837 270
837 288
0 1 20 0 0 4224 0 0 17 57 0 2
613 270
702 270
2 1 18 0 0 0 0 44 18 0 0 2
297 270
360 270
1 0 21 0 0 4096 0 19 0 0 61 2
522 117
522 135
1 2 2 0 0 128 0 40 23 0 0 5
414 333
414 354
406 354
406 329
202 329
1 0 2 0 0 0 0 20 0 0 58 2
504 354
504 354
1 0 2 0 0 128 0 39 0 0 58 3
837 324
837 345
504 345
2 3 20 0 0 0 0 41 22 0 0 3
612 297
613 297
613 226
3 0 2 0 0 0 0 21 0 0 0 2
504 288
504 360
0 2 22 0 0 4096 0 0 22 60 0 2
521 208
590 208
1 1 22 0 0 8320 0 21 42 0 0 4
504 252
521 252
521 180
522 180
0 1 21 0 0 8192 0 0 22 62 0 4
522 136
522 135
613 135
613 190
2 2 21 0 0 8320 0 43 42 0 0 4
414 144
414 136
522 136
522 144
1 1 23 0 0 4224 0 23 44 0 0 4
202 319
253 319
253 270
261 270
0
0
2073 0 1
0
0
0
0 0 0
0
0 0 0
100 1 0.01 1e+008
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
2 0 0 0
2 Rf
1000 10000 9000
3 Rf1
1e+006 1e+007 9e+006
5 -1 10 10 10 0 10 10 0
1444834 1210432 100 100 0 0
0 0 0 0
0 71 161 141
0 66
0 66
1247 66
1247 396
0 0
0 0 0 0 0 0
12401 0
4 0.3 10
1
837 280
0 17 0 0 2	0 50 0 0
2818758 8813120 100 100 0 0
77 66 977 426
1025 79 2049 595
977 66
77 66
977 94
977 401
0 0
0.005 0 1.78182e-008 -1.80727e-008 0.005 0.005
28921 0
4 0.001 10
1
837 290
0 17 0 0 2	39 0 0 0
5046462 4421696 100 100 0 0
77 66 987 426
1025 595 2049 1111
715 66
715 66
987 122
987 235
0 0
103587 103587 41.4815 3.7037 1e+008 1e+008
12530 0
4 3e+007 5e+007
11
819 270
0 17 0 0 1	0 50 0 0
819 270
0 17 0 0 1	0 50 0 0
819 270
0 17 0 0 1	0 50 0 0
819 270
0 17 0 0 1	0 50 0 0
819 270
0 17 0 0 1	0 50 0 0
811 972
0 3 0 0 1	0 8 0 0
802 625
0 10 0 0 1	0 29 0 0
802 625
0 10 0 0 1	0 29 0 0
802 625
0 10 0 0 1	0 29 0 0
802 625
0 10 0 0 1	0 29 0 0
802 625
0 10 0 0 1	0 29 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
